* E:\2-1\EEE 210\Schematics\main.sch

* Schematics Version 9.2
* Mon Jun 06 20:51:10 2016



** Analysis setup **
.tran 1ns 5m 0 1u
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "main.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
